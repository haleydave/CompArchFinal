module imem(CLK, instr, ADD);

input CLK;
output [15:0] instr;
input [2:0] ADD; 

//input reg and stuff to read from assembled file after I actually figure out assembler


endmodule